library ieee;
use ieee.std_logic_1164.all;


entity subbyte is
	port (
		clk		: in  std_logic;
		input	: in  std_logic_vector(7 downto 0);
		output	: out std_logic_vector(7 downto 0)
	);
end entity;


architecture subbyte_arch of subbyte is
begin
	process (clk)
	begin
		if rising_edge(clk) then
			case input is
				when X"00" => output <= X"63";
				when X"01" => output <= X"7c";
				when X"02" => output <= X"77";
				when X"03" => output <= X"7b";
				when X"04" => output <= X"f2";
				when X"05" => output <= X"6b";
				when X"06" => output <= X"6f";
				when X"07" => output <= X"c5";
				when X"08" => output <= X"30";
				when X"09" => output <= X"01";
				when X"0a" => output <= X"67";
				when X"0b" => output <= X"2b";
				when X"0c" => output <= X"fe";
				when X"0d" => output <= X"d7";
				when X"0e" => output <= X"ab";
				when X"0f" => output <= X"76";
				when X"10" => output <= X"ca";
				when X"11" => output <= X"82";
				when X"12" => output <= X"c9";
				when X"13" => output <= X"7d";
				when X"14" => output <= X"fa";
				when X"15" => output <= X"59";
				when X"16" => output <= X"47";
				when X"17" => output <= X"f0";
				when X"18" => output <= X"ad";
				when X"19" => output <= X"d4";
				when X"1a" => output <= X"a2";
				when X"1b" => output <= X"af";
				when X"1c" => output <= X"9c";
				when X"1d" => output <= X"a4";
				when X"1e" => output <= X"72";
				when X"1f" => output <= X"c0";
				when X"20" => output <= X"b7";
				when X"21" => output <= X"fd";
				when X"22" => output <= X"93";
				when X"23" => output <= X"26";
				when X"24" => output <= X"36";
				when X"25" => output <= X"3f";
				when X"26" => output <= X"f7";
				when X"27" => output <= X"cc";
				when X"28" => output <= X"34";
				when X"29" => output <= X"a5";
				when X"2a" => output <= X"e5";
				when X"2b" => output <= X"f1";
				when X"2c" => output <= X"71";
				when X"2d" => output <= X"d8";
				when X"2e" => output <= X"31";
				when X"2f" => output <= X"15";
				when X"30" => output <= X"04";
				when X"31" => output <= X"c7";
				when X"32" => output <= X"23";
				when X"33" => output <= X"c3";
				when X"34" => output <= X"18";
				when X"35" => output <= X"96";
				when X"36" => output <= X"05";
				when X"37" => output <= X"9a";
				when X"38" => output <= X"07";
				when X"39" => output <= X"12";
				when X"3a" => output <= X"80";
				when X"3b" => output <= X"e2";
				when X"3c" => output <= X"eb";
				when X"3d" => output <= X"27";
				when X"3e" => output <= X"b2";
				when X"3f" => output <= X"75";
				when X"40" => output <= X"09";
				when X"41" => output <= X"83";
				when X"42" => output <= X"2c";
				when X"43" => output <= X"1a";
				when X"44" => output <= X"1b";
				when X"45" => output <= X"6e";
				when X"46" => output <= X"5a";
				when X"47" => output <= X"a0";
				when X"48" => output <= X"52";
				when X"49" => output <= X"3b";
				when X"4a" => output <= X"d6";
				when X"4b" => output <= X"b3";
				when X"4c" => output <= X"29";
				when X"4d" => output <= X"e3";
				when X"4e" => output <= X"2f";
				when X"4f" => output <= X"84";
				when X"50" => output <= X"53";
				when X"51" => output <= X"d1";
				when X"52" => output <= X"00";
				when X"53" => output <= X"ed";
				when X"54" => output <= X"20";
				when X"55" => output <= X"fc";
				when X"56" => output <= X"b1";
				when X"57" => output <= X"5b";
				when X"58" => output <= X"6a";
				when X"59" => output <= X"cb";
				when X"5a" => output <= X"be";
				when X"5b" => output <= X"39";
				when X"5c" => output <= X"4a";
				when X"5d" => output <= X"4c";
				when X"5e" => output <= X"58";
				when X"5f" => output <= X"cf";
				when X"60" => output <= X"d0";
				when X"61" => output <= X"ef";
				when X"62" => output <= X"aa";
				when X"63" => output <= X"fb";
				when X"64" => output <= X"43";
				when X"65" => output <= X"4d";
				when X"66" => output <= X"33";
				when X"67" => output <= X"85";
				when X"68" => output <= X"45";
				when X"69" => output <= X"f9";
				when X"6a" => output <= X"02";
				when X"6b" => output <= X"7f";
				when X"6c" => output <= X"50";
				when X"6d" => output <= X"3c";
				when X"6e" => output <= X"9f";
				when X"6f" => output <= X"a8";
				when X"70" => output <= X"51";
				when X"71" => output <= X"a3";
				when X"72" => output <= X"40";
				when X"73" => output <= X"8f";
				when X"74" => output <= X"92";
				when X"75" => output <= X"9d";
				when X"76" => output <= X"38";
				when X"77" => output <= X"f5";
				when X"78" => output <= X"bc";
				when X"79" => output <= X"b6";
				when X"7a" => output <= X"da";
				when X"7b" => output <= X"21";
				when X"7c" => output <= X"10";
				when X"7d" => output <= X"ff";
				when X"7e" => output <= X"f3";
				when X"7f" => output <= X"d2";
				when X"80" => output <= X"cd";
				when X"81" => output <= X"0c";
				when X"82" => output <= X"13";
				when X"83" => output <= X"ec";
				when X"84" => output <= X"5f";
				when X"85" => output <= X"97";
				when X"86" => output <= X"44";
				when X"87" => output <= X"17";
				when X"88" => output <= X"c4";
				when X"89" => output <= X"a7";
				when X"8a" => output <= X"7e";
				when X"8b" => output <= X"3d";
				when X"8c" => output <= X"64";
				when X"8d" => output <= X"5d";
				when X"8e" => output <= X"19";
				when X"8f" => output <= X"73";
				when X"90" => output <= X"60";
				when X"91" => output <= X"81";
				when X"92" => output <= X"4f";
				when X"93" => output <= X"dc";
				when X"94" => output <= X"22";
				when X"95" => output <= X"2a";
				when X"96" => output <= X"90";
				when X"97" => output <= X"88";
				when X"98" => output <= X"46";
				when X"99" => output <= X"ee";
				when X"9a" => output <= X"b8";
				when X"9b" => output <= X"14";
				when X"9c" => output <= X"de";
				when X"9d" => output <= X"5e";
				when X"9e" => output <= X"0b";
				when X"9f" => output <= X"db";
				when X"a0" => output <= X"e0";
				when X"a1" => output <= X"32";
				when X"a2" => output <= X"3a";
				when X"a3" => output <= X"0a";
				when X"a4" => output <= X"49";
				when X"a5" => output <= X"06";
				when X"a6" => output <= X"24";
				when X"a7" => output <= X"5c";
				when X"a8" => output <= X"c2";
				when X"a9" => output <= X"d3";
				when X"aa" => output <= X"ac";
				when X"ab" => output <= X"62";
				when X"ac" => output <= X"91";
				when X"ad" => output <= X"95";
				when X"ae" => output <= X"e4";
				when X"af" => output <= X"79";
				when X"b0" => output <= X"e7";
				when X"b1" => output <= X"c8";
				when X"b2" => output <= X"37";
				when X"b3" => output <= X"6d";
				when X"b4" => output <= X"8d";
				when X"b5" => output <= X"d5";
				when X"b6" => output <= X"4e";
				when X"b7" => output <= X"a9";
				when X"b8" => output <= X"6c";
				when X"b9" => output <= X"56";
				when X"ba" => output <= X"f4";
				when X"bb" => output <= X"ea";
				when X"bc" => output <= X"65";
				when X"bd" => output <= X"7a";
				when X"be" => output <= X"ae";
				when X"bf" => output <= X"08";
				when X"c0" => output <= X"ba";
				when X"c1" => output <= X"78";
				when X"c2" => output <= X"25";
				when X"c3" => output <= X"2e";
				when X"c4" => output <= X"1c";
				when X"c5" => output <= X"a6";
				when X"c6" => output <= X"b4";
				when X"c7" => output <= X"c6";
				when X"c8" => output <= X"e8";
				when X"c9" => output <= X"dd";
				when X"ca" => output <= X"74";
				when X"cb" => output <= X"1f";
				when X"cc" => output <= X"4b";
				when X"cd" => output <= X"bd";
				when X"ce" => output <= X"8b";
				when X"cf" => output <= X"8a";
				when X"d0" => output <= X"70";
				when X"d1" => output <= X"3e";
				when X"d2" => output <= X"b5";
				when X"d3" => output <= X"66";
				when X"d4" => output <= X"48";
				when X"d5" => output <= X"03";
				when X"d6" => output <= X"f6";
				when X"d7" => output <= X"0e";
				when X"d8" => output <= X"61";
				when X"d9" => output <= X"35";
				when X"da" => output <= X"57";
				when X"db" => output <= X"b9";
				when X"dc" => output <= X"86";
				when X"dd" => output <= X"c1";
				when X"de" => output <= X"1d";
				when X"df" => output <= X"9e";
				when X"e0" => output <= X"e1";
				when X"e1" => output <= X"f8";
				when X"e2" => output <= X"98";
				when X"e3" => output <= X"11";
				when X"e4" => output <= X"69";
				when X"e5" => output <= X"d9";
				when X"e6" => output <= X"8e";
				when X"e7" => output <= X"94";
				when X"e8" => output <= X"9b";
				when X"e9" => output <= X"1e";
				when X"ea" => output <= X"87";
				when X"eb" => output <= X"e9";
				when X"ec" => output <= X"ce";
				when X"ed" => output <= X"55";
				when X"ee" => output <= X"28";
				when X"ef" => output <= X"df";
				when X"f0" => output <= X"8c";
				when X"f1" => output <= X"a1";
				when X"f2" => output <= X"89";
				when X"f3" => output <= X"0d";
				when X"f4" => output <= X"bf";
				when X"f5" => output <= X"e6";
				when X"f6" => output <= X"42";
				when X"f7" => output <= X"68";
				when X"f8" => output <= X"41";
				when X"f9" => output <= X"99";
				when X"fa" => output <= X"2d";
				when X"fb" => output <= X"0f";
				when X"fc" => output <= X"b0";
				when X"fd" => output <= X"54";
				when X"fe" => output <= X"bb";
				when X"ff" => output <= X"16";
				when others => output <= X"FF";
			end case;
		end if;
	end process;
end architecture;
